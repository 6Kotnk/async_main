`timescale 1ns / 1ps

module top_wraper();
/*
(* DONT_TOUCH = "yes" *)
module top_wraper(

  output [7:0] JA,

  input btnC,
  
  input clk
);

fib_tp_top TOP
(
//---------CTRL-----------------------
  .clk                        (clk),
  .btnC                       (btnC),
//---------IO-------------------------
  .JA                         (JA)
//------------------------------------
);
*/
endmodule