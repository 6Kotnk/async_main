package link_pkg;
parameter RAIL_NUM = 2;

typedef logic [RAIL_NUM-1:0] multi_rail_bit;

endpackage