`timescale 1ns / 1ps

module top_wraper(
  input clk
);


endmodule